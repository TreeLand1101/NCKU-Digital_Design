// 
// Designer: P76124265
//

module Max_Heapify(Array, Size, index, enble, done);

endmodule

module Build_Queue(Array, Size, enble, done);

endmodule

module Extract_Max(Array, Size, enble, done);

endmodule

module Increase_Value(Array, Size, index, value, enble, done);

endmodule

module Insert_Data(Array, Size, value, enble, done);

endmodule