module shiftRows_tb;

reg [127:0] in;
wire [127:0] out;	


shiftRows m (in,out);


initial begin
	$monitor("input= %H , output= %h, ans = d4bf5d30e0b452aeb84111f11e2798e5",in,out);
	in = 128'hd42711aee0bf98f1b8b45de51e415230;
end
endmodule